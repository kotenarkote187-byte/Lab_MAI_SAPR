`timescale 1ns/1ps

module apb_slave (
    // ????????? APB ????
    input  logic        PCLK,      // ???????? ??????
    input  logic        PRESETn,   // ????? (???????? ?????? ???????)
    input  logic        PSEL,      // ????? ???????? ??????????
    input  logic        PENABLE,   // ?????????? ????????
    input  logic        PWRITE,   // ??????????? ???????? (1-??????, 0-??????)
    input  logic [31:0] PADDR,    // ????? ????
    input  logic [31:0] PWDATA,   // ?????? ??? ??????
    output logic [31:0] PRDATA,   // ?????? ??? ??????
    output logic        PREADY,   // ?????????? ????????
    output logic        PSLVERR   // ?????? ????????
);

    // ?????????? ???????? ??? ???????? ?????? (16 ????????? ?? 32 ????)
    logic [31:0] registers [0:15];
    
    // ??????? ?????????? ?????? ?????? ? ?? ?????????? ??????
    assign PREADY = 1'b1;   // ?????? ????? ? ???????????
    assign PSLVERR = 1'b0;  // ?????? ???????????

    // ?????? ?????? ? ???????? (??????????)
    always_ff @(posedge PCLK or negedge PRESETn) begin
        if (!PRESETn) begin
            // ????? ???? ????????? ? 0
            foreach(registers[i]) begin
                registers[i] <= 32'd0;
            end
            $display("");
            $display("================================================");
            $display("APB ??????? ??????????: ????? ????????");
            $display("??? ???????? ???????????????? ? 0x00000000");
            $display("================================================");
            $display("");
        end else if (PSEL && PENABLE && PWRITE) begin
            // ???????? ??????: PSEL=1, PENABLE=1, PWRITE=1
            if (PADDR[31:4] == 28'h0) begin
                // ?????? ? ??????? (?????? 0x0 - 0xF)
                registers[PADDR[3:0]] <= PWDATA;
                $display("");
                $display("------------------------------------------------");
                $display("APB ??????? ??????????: ???????? ??????");
                $display("------------------------------------------------");
                $display("???????[0x%01h] = 0x%08h", PADDR[3:0], PWDATA);
                $display("?????????? ????????: 0x%08h", registers[PADDR[3:0]]);
                $display("?????? ??????? ?????????");
                $display("------------------------------------------------");
                $display("");
            end else begin
                // ???????????? ????? ??? ??????
                $display("APB ??????? ??????????: ???????? ????? ?????? 0x%08h", PADDR);
            end
        end
    end

    // ?????? ?????? ?? ????????? - ?????????????? ?????? ??? ???????????? ??????
    always_comb begin
        PRDATA = 32'd0;  // ???????? ?? ?????????
        if (PSEL && !PWRITE) begin
            // ???????? ??????: PSEL=1, PWRITE=0
            if (PADDR[31:4] == 28'h0) begin
                // ?????? ?? ???????? (?????? 0x0 - 0xF)
                PRDATA = registers[PADDR[3:0]];
                $display("");
                $display("------------------------------------------------");
                $display("APB ??????? ??????????: ???????? ?????? - ??????????????");
                $display("------------------------------------------------");
                $display("?????? ????????[0x%01h]", PADDR[3:0]);
                $display("?????? ??? ??????: 0x%08h", registers[PADDR[3:0]]);
                $display("PRDATA ?????????? ?: 0x%08h", PRDATA);
                $display("?????? ??? ?????? ?????? ??????????");
                $display("------------------------------------------------");
                $display("");
            end else begin
                // ???????????? ????? ??? ?????? - ?????????? ???????? ????????
                PRDATA = 32'hDEADBEEF;
                $display("APB ??????? ??????????: ???????? ????? ?????? 0x%08h, ????????? 0xDEADBEEF", PADDR);
            end
        end
    end

    // ??????? ??? ??????? - ?????? ???? ?????????
    function void print_all_registers();
        begin
            $display("");
            $display("================================================");
            $display("APB ??????? ??????????: ???? ?????????");
            $display("================================================");
            for (int i = 0; i < 16; i++) begin
                $display("???????[0x%01h] = 0x%08h", i, registers[i]);
            end
            $display("================================================");
            $display("");
        end
    endfunction

endmodule