`timescale 1ns/1ps

module Testbench;

    // ???????? ?????? ? ?????
    logic clk;
    logic rst_n;
    
    // APB ??????? (Advanced Peripheral Bus)
    logic        PSEL;      // ????? ???????? ??????????
    logic        PENABLE;   // ?????????? ????????
    logic        PWRITE;   // ??????????? ???????? (1-??????, 0-??????)
    logic [31:0] PADDR;    // ????? ????
    logic [31:0] PWDATA;   // ?????? ??? ??????
    logic [31:0] PRDATA;   // ?????? ??? ??????
    logic        PREADY;   // ?????????? ????????
    logic        PSLVERR;  // ?????? ????????
    
    // ????????? ????????? ???????
    initial begin
        clk = 0;
        $display("?????? ????????? ????????? ???????...");
        forever #5 clk = ~clk;  // ?????? 10 ?? (??????? 100 ???)
    end
    
    // ????????? ??????? ??????
    initial begin
        rst_n = 0;  // ???????? ?????? ??????? ??????
        $display("????? ???????????");
        #20 rst_n = 1;  // ?????? ?????? ????? 20 ??
        $display("????? ???? ? ?????? ??????? %0t", $time);
    end
    
    // ????????? ??????? APB (??????? ??????????)
    apb_master master_inst (
        .PCLK(clk),
        .PRESETn(rst_n),
        .PSEL(PSEL),
        .PENABLE(PENABLE),
        .PWRITE(PWRITE),
        .PADDR(PADDR),
        .PWDATA(PWDATA),
        .PRDATA(PRDATA),
        .PREADY(PREADY),
        .PSLVERR(PSLVERR)
    );
    
    // ????????? ?????? APB (??????? ??????????)
    apb_slave slave_inst (
        .PCLK(clk),
        .PRESETn(rst_n),
        .PSEL(PSEL),
        .PENABLE(PENABLE),
        .PWRITE(PWRITE),
        .PADDR(PADDR),
        .PWDATA(PWDATA),
        .PRDATA(PRDATA),
        .PREADY(PREADY),
        .PSLVERR(PSLVERR)
    );
    
    // ???????? ???????? ????????
    initial begin
        logic [31:0] read_data;  // ?????????? ??? ???????? ??????????? ??????
        
        // ???????? ?????????? ??????
        #30;
        $display("");
        $display("************************************************");
        $display("???????????? APB ??????? ??????");
        $display("************************************************");
        $display("");
        
        // 1. ?????? ???????? 2 ?? ?????? 0x0
        $display("???? 1: ?????? ???????? 2 ?? ?????? 0x0");
        master_inst.apb_write(32'h00000000, 32'h00000002);
        #50;  // ???????? 50 ??
        
        // 2. ?????? ???? ?? ?????? 0x4
        $display("???? 2: ?????? ???? ?? ?????? 0x4");
        master_inst.apb_write(32'h00000004, 32'h15122024);  // 15.12.2024
        #50;
        
        // 3. ?????? ??????? ?? ?????? 0x8
        $display("???? 3: ?????? ??????? ?? ?????? 0x8");
        master_inst.apb_write(32'h00000008, 32'h4D49524F); // MIRO ? ASCII
        #50;

        // 4. ?????? ????? ?? ?????? 0xC
        $display("???? 4: ?????? ????? ?? ?????? 0xC");
        master_inst.apb_write(32'h0000000C, 32'h45474F52); // EGOR ? ASCII
        #50;
        
        // ?????? ???? ????????? ?????? ??? ????????
        slave_inst.print_all_registers();
        
        // ???? ??????????? - ?????? ?????????? ??????
        $display("");
        $display("************************************************");
        $display("???? ????????: ?????? ???? ?????????? ????????");
        $display("************************************************");
        $display("");
        
        // ?????? ?????? 0x0
        $display("?????? ?????? 0x0");
        master_inst.apb_read(32'h00000000, read_data);
        $display("????????: ????????? ? ?????? 0x0 = 0x%08h (?????????: 0x00000002)", read_data);
        if (read_data == 32'h00000002) 
            $display("?????: ?????? ????????????? ?????????? ????????!");
        else 
            $display("??????: ?????????????? ??????!");
        #20;
        
        // ?????? ?????? 0x4
        $display("?????? ?????? 0x4");
        master_inst.apb_read(32'h00000004, read_data);
        $display("????????: ????????? ? ?????? 0x4 = 0x%08h (?????????: 0x15122024)", read_data);
        if (read_data == 32'h15122024) 
            $display("?????: ?????? ????????????? ?????????? ????????!");
        else 
            $display("??????: ?????????????? ??????!");
        #20;
        
        // ?????? ?????? 0x8
        $display("?????? ?????? 0x8");
        master_inst.apb_read(32'h00000008, read_data);
        $display("????????: ????????? ? ?????? 0x8 = 0x%08h (?????????: 0x4D49524F)", read_data);
        if (read_data == 32'h4D49524F) 
            $display("?????: ?????? ????????????? ?????????? ????????!");
        else 
            $display("??????: ?????????????? ??????!");
        #20;
        
        // ?????? ?????? 0xC
        $display("?????? ?????? 0xC");
        master_inst.apb_read(32'h0000000C, read_data);
        $display("????????: ????????? ? ?????? 0xC = 0x%08h (?????????: 0x45474F52)", read_data);
        if (read_data == 32'h45474F52) 
            $display("?????: ?????? ????????????? ?????????? ????????!");
        else 
            $display("??????: ?????????????? ??????!");
        #20;
        
        // ????????? ?????
        $display("");
        $display("************************************************");
        $display("???????????? APB ??????? ?????????");
        $display("************************************************");
        $display("????: ??? ???????? ?????????");
        $display("????? ?????????: %0t ??", $time);
        $display("************************************************");
        $display("");
        
        #50;
        $finish;  // ?????????? ?????????
    end
    
    // ?????????? ???? APB ? ???????? ???????
    initial begin
        $monitor("?????: %0t | APB_????: PSEL=%b PENABLE=%b PWRITE=%b PADDR=0x%08h PWDATA=0x%08h PRDATA=0x%08h PREADY=%b", 
                 $time, PSEL, PENABLE, PWRITE, PADDR, PWDATA, PRDATA, PREADY);
    end

    // ????-??? ??? ???????????? (?? ?????? ????????? ?????????)
    initial begin
        #2000;  // ????-??? 2000 ??
        $display("");
        $display("????-???: ????????? ?????? ??????? ????? ???????, ?????????????? ??????????");
        $display("");
        $finish;
    end

endmodule